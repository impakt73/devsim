`ifndef PKG_COMMON
`define PKG_COMMON

package common;

typedef enum
{
    mem_req_size_byte,
    mem_req_size_half,
    mem_req_size_word
} mem_req_size;

endpackage

`endif